.subckt inv in out VDD VSS
Mp out in VDD VDD p_18 w=wp l=len
Mn out in VSS VSS n_18 w=wn l=len
.ends