.subckt mux_arr a0 a1 a2 a3 a4 a5 a6 a7 a8 a9 a10 a11 a12 a13 a14 a15
+ b0 b1 b2 b3 b4 b5 b6 b7 b8 b9 b10 b11 b12 b13 b14 b15 S
+ out0 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15 VDD VSS
Xmux0 a0 b0 S out0 VDD VSS mux m=1
Xmux1 a1 b1 S out1 VDD VSS mux m=1
Xmux2 a2 b2 S out2 VDD VSS mux m=1
Xmux3 a3 b3 S out3 VDD VSS mux m=1
Xmux4 a4 b4 S out4 VDD VSS mux m=1
Xmux5 a5 b5 S out5 VDD VSS mux m=1
Xmux6 a6 b6 S out6 VDD VSS mux m=1
Xmux7 a7 b7 S out7 VDD VSS mux m=1
Xmux8 a8 b8 S out8 VDD VSS mux m=1
Xmux9 a9 b9 S out9 VDD VSS mux m=1
Xmux10 a10 b10 S out10 VDD VSS mux m=1
Xmux11 a11 b11 S out11 VDD VSS mux m=1
Xmux12 a12 b12 S out12 VDD VSS mux m=1
Xmux13 a13 b13 S out13 VDD VSS mux m=1
Xmux14 a14 b14 S out14 VDD VSS mux m=1
Xmux15 a15 b15 S out15 VDD VSS mux m=1
.ends