.subckt ff_arr clk in0 in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15
+ out0 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15
+ outb0 outb1 outb2 outb3 outb4 outb5 outb6 outb7 outb8 outb9 outb10 outb11 outb12 outb13 outb14 outb15 VDD VSS
Xff0 clk in0 out0 outb0 VDD VSS ff m=1
Xff1 clk in1 out1 outb1 VDD VSS ff m=1
Xff2 clk in2 out2 outb2 VDD VSS ff m=1
Xff3 clk in3 out3 outb3 VDD VSS ff m=1
Xff4 clk in4 out4 outb4 VDD VSS ff m=1
Xff5 clk in5 out5 outb5 VDD VSS ff m=1
Xff6 clk in6 out6 outb6 VDD VSS ff m=1
Xff7 clk in7 out7 outb7 VDD VSS ff m=1
Xff8 clk in8 out8 outb8 VDD VSS ff m=1
Xff9 clk in9 out9 outb9 VDD VSS ff m=1
Xff10 clk in10 out10 outb10 VDD VSS ff m=1
Xff11 clk in11 out11 outb11 VDD VSS ff m=1
Xff12 clk in12 out12 outb12 VDD VSS ff m=1
Xff13 clk in13 out13 outb13 VDD VSS ff m=1
Xff14 clk in14 out14 outb14 VDD VSS ff m=1
Xff15 clk in15 out15 outb15 VDD VSS ff m=1
.ends
