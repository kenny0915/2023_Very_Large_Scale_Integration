.subckt inv_arr in0 in1 in2 in3 in4 in5 in6 in7 in8 in9 in10 in11 in12 in13 in14 in15
+ out0 out1 out2 out3 out4 out5 out6 out7 out8 out9 out10 out11 out12 out13 out14 out15 VDD VSS
Xinv0 in0 out0 VDD VSS inv m=1
Xinv1 in1 out1 VDD VSS inv m=1 
Xinv2 in2 out2 VDD VSS inv m=1 
Xinv3 in3 out3 VDD VSS inv m=1
Xinv4 in4 out4 VDD VSS inv m=1 
Xinv5 in5 out5 VDD VSS inv m=1 
Xinv6 in6 out6 VDD VSS inv m=1 
Xinv7 in7 out7 VDD VSS inv m=1 
Xinv8 in8 out8 VDD VSS inv m=1
Xinv9 in9 out9 VDD VSS inv m=1 
Xinv10 in10 out10 VDD VSS inv m=1
Xinv11 in11 out11 VDD VSS inv m=1
Xinv12 in12 out12 VDD VSS inv m=1
Xinv13 in13 out13 VDD VSS inv m=1
Xinv14 in14 out14 VDD VSS inv m=1
Xinv15 in15 out15 VDD VSS inv m=1
.ends